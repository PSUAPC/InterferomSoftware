LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;

entity IntegratorCLPD_tb is
end entity IntegratorCLPD_tb;
architecture RTL of IntegratorCLPD_tb is
--Signals and components go here
component IntegratorCLPD is
port(
 -- comparison variables
 pulse : in std_logic;
 latch : in std_logic;
 dataIn : in std_logic;
 output : out std_logic;
 loaded : out std_logic;
 
 -- count variables
 fvcIn : in std_logic;
 wordSelect : in std_logic;
 dataOut : out std_logic_vector(15 downto 0)
 );
end component IntegratorCLPD;

signal pulse: std_logic;
signal latch: std_logic;
signal dataIn : std_logic;
signal output : std_logic;
signal loaded : std_logic;

signal fvcIn: std_logic;
signal wordSelect: std_logic;
signal dataOut : std_logic_vector(15 downto 0);

begin

	DUT: IntegratorCLPD port map( pulse => pulse, latch => latch, dataIn => dataIn, output => output, 
									loaded => loaded, fvcIn => fvcIn, wordSelect => wordSelect, dataOut => dataOut);
	
	process
	begin
	-- set the signals to null
	pulse <= '0';
	latch <= '0';
	dataIn <= '0';
	fvcIn <= '0';
	wordSelect <= '0';
									
	-- lets shift in a number
	for i in 0 to 28 loop
	  latch <= '1';
	  wait for 10 ns;
	  latch <= '0';
	  wait for 10 ns;
	end loop;
	
	dataIn <= '1';
	
	for i in 0 to 2 loop
		latch <= '1';
	  wait for 10 ns;
	  latch <= '0';
	  wait for 10 ns;  
	end loop;
	
	-- reload again for testing
	dataIn <= '0';
	for i in 0 to 28 loop
	  latch <= '1';
	  wait for 10 ns;
	  latch <= '0';
	  wait for 10 ns;
	end loop;
	
	dataIn <= '1';
	
	for i in 0 to 2 loop
		latch <= '1';
	  wait for 10 ns;
	  latch <= '0';
	  wait for 10 ns;  
	end loop;
	
		-- reload again for testing
	dataIn <= '0';
	for i in 0 to 28 loop
	  latch <= '1';
	  wait for 10 ns;
	  latch <= '0';
	  wait for 10 ns;
	end loop;
	
	dataIn <= '1';
	
	for i in 0 to 2 loop
		latch <= '1';
	  wait for 10 ns;
	  latch <= '0';
	  wait for 10 ns;  
	end loop;
	
	-- now, lets start pulsing
  for i in 0 to 20 loop
	  pulse <= '1';
	  wait for 10 ns;
	  pulse <= '0';
	  wait for 10 ns;
	end loop;
	
	fvcIn <= '1';
	wait for 10 ns;
	fvcIn <= '0';
	wait for 10 ns;
	
	pulse <= '1';
	wait for 10 ns;
	pulse <= '0';
	wait for 10 ns;
	
  fvcIn <= '1';
	wait for 10 ns;
	fvcIn <= '0';
	wait for 10 ns;
	
	for i in 0 to 4 loop
	  pulse <= '1';
	  wait for 10 ns;
	  pulse <= '0';
	  wait for 10 ns;
	end loop;
	
		pulse <= '1';
		fvcIn <= '1';
	  wait for 10 ns;
	  pulse <= '0';
	  fvcIn <= '0';
	  wait for 10 ns;
	
			pulse <= '1';
		fvcIn <= '1';
	  wait for 10 ns;
	  pulse <= '0';
	  fvcIn <= '0';
	  wait for 10 ns;
	  
	  		pulse <= '1';
		fvcIn <= '1';
	  wait for 10 ns;
	  pulse <= '0';
	  fvcIn <= '0';
	  wait for 10 ns;
	  
		for i in 0 to 12 loop
	   pulse <= '1';
	   wait for 10 ns;
	   pulse <= '0';
	   wait for 10 ns;
	  end loop;
	  
	  			pulse <= '1';
		fvcIn <= '1';
	  wait for 10 ns;
	  pulse <= '0';
	  fvcIn <= '0';
	  wait for 10 ns;
	  
	  		pulse <= '1';
		fvcIn <= '1';
	  wait for 10 ns;
	  pulse <= '0';
	  fvcIn <= '0';
	  wait for 10 ns;

	  		pulse <= '1';
		fvcIn <= '1';
	  wait for 10 ns;
	  pulse <= '0';
	  fvcIn <= '0';
	  wait for 10 ns;
	  
	  	  		pulse <= '1';
		fvcIn <= '1';
	  wait for 10 ns;
	  pulse <= '0';
	  fvcIn <= '0';
	  wait for 10 ns;
	  	  
		for i in 0 to 6 loop
	   pulse <= '1';
	   wait for 10 ns;
	   pulse <= '0';
	   wait for 10 ns;
	  end loop;
	  
	  	  		pulse <= '1';
		fvcIn <= '1';
	  wait for 10 ns;
	  pulse <= '0';
	  fvcIn <= '0';
	  wait for 10 ns;
	  
	  	  		pulse <= '1';
		fvcIn <= '1';
	  wait for 10 ns;
	  pulse <= '0';
	  fvcIn <= '0';
	  wait for 10 ns;
	  
	  		for i in 0 to 2 loop
	   pulse <= '1';
	   wait for 10 ns;
	   pulse <= '0';
	   wait for 10 ns;
	  end loop;
	  
	  pulse <= '1';
		latch <= '1';
	  wait for 10 ns;
	  pulse <= '0';
	  latch <= '0';
	  wait for 10 ns;
	
		  		for i in 0 to 12 loop
	   pulse <= '1';
	   wait for 10 ns;
	   pulse <= '0';
	   wait for 10 ns;
	  end loop;
	  
	wait;
	end process;

end architecture RTL;