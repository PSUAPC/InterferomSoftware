LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;

entity FlagRegister is
generic (N : integer);
port(
 -- comparison variables
 clk : in std_logic;
 reset : in std_logic;
 regIn : in std_logic_vector(N-1 downto 0);
 
 regOut : out std_logic_vector(N-1 downto 0)
 );
end entity FlagRegister;

architecture RTL of FlagRegister is

signal reg : std_logic_vector(N-1 downto 0) :=  (others =>'0');

begin

	-- define the flag or process
	process( clk, reset )

	begin
		-- synchronous reset
		if(rising_edge(clk) ) then
			if( reset = '1') then
				reg <= (others =>'0');
			else 
				reg <= reg OR regIn;
			end if;
		end if;
	end process;

	-- link the output
	regOut <= reg;

end architecture RTL;